package axis2nas_pkg is
	constant AXI_BUS_BIT_WIDTH : integer := 32;
	constant NAS_CONFIG_BUS_BIT_WIDTH : integer := 16;
end package axis2nas_pkg;

package body axis2nas_pkg is
end package body axis2nas_pkg;
