--///////////////////////////////////////////////////////////////////////////////
--//                                                                           //
--//    Copyright © 2016  Angel Francisco Jimenez-Fernandez                    //
--//                                                                           //
--//    This file is part of OpenNAS.                                          //
--//                                                                           //
--//    OpenNAS is free software: you can redistribute it and/or modify        //
--//    it under the terms of the GNU General Public License as published by   //
--//    the Free Software Foundation, either version 3 of the License, or      //
--//    (at your option) any later version.                                    //
--//                                                                           //
--//    OpenNAS is distributed in the hope that it will be useful,             //
--//    but WITHOUT ANY WARRANTY; without even the implied warranty of         //
--//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.See the            //
--//    GNU General Public License for more details.                           //
--//                                                                           //
--//    You should have received a copy of the GNU General Public License      //
--//    along with OpenNAS. If not, see <http://www.gnu.org/licenses/>.        //
--//                                                                           //
--///////////////////////////////////////////////////////////////////////////////

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;           -- @suppress "Deprecated package"
use ieee.std_logic_unsigned.all;        -- @suppress "Deprecated package"
use work.OpenNas_top_pkg.all;
use ieee.numeric_std.all;

entity CFBank_2or_8CH is
	generic(
		CONFIG_ADDRESS : integer := 16#0000#;
		CONFIG_OFFSET  : integer := 35  -- Don't change this value
	);
	Port(
		clock       : in  std_logic;
		rst         : in  std_logic;
		--Config Bus
		config_data : in  std_logic_vector(CONFIG_BUS_BIT_WIDTH - 1 downto 0);
		config_addr : in  std_logic_vector(CONFIG_BUS_BIT_WIDTH - 1 downto 0);
		config_wren : in  std_logic;
		--Output
		spikes_in   : in  std_logic_vector(1 downto 0);
		spikes_out  : out std_logic_vector(15 downto 0)
	);
end CFBank_2or_8CH;

architecture CFBank_arq of CFBank_2or_8CH is

	signal not_rst      : std_logic;
	signal lpf_spikes_0 : std_logic_vector(1 downto 0);
	signal lpf_spikes_1 : std_logic_vector(1 downto 0);
	signal lpf_spikes_2 : std_logic_vector(1 downto 0);
	signal lpf_spikes_3 : std_logic_vector(1 downto 0);
	signal lpf_spikes_4 : std_logic_vector(1 downto 0);
	signal lpf_spikes_5 : std_logic_vector(1 downto 0);
	signal lpf_spikes_6 : std_logic_vector(1 downto 0);
	signal lpf_spikes_7 : std_logic_vector(1 downto 0);
	signal lpf_spikes_8 : std_logic_vector(1 downto 0); -- @suppress "signal lpf_spikes_8 is never read"

	-- Configurable signals
	type register_bank is array (0 to CONFIG_OFFSET) of std_logic_vector(CONFIG_BUS_BIT_WIDTH - 1 downto 0);
	signal config_mem : register_bank;

begin

	not_rst <= not rst;

	U_Config_registers : process(clock, not_rst)
	begin
		if (not_rst = '0') then         -- In reset mode the parameter are the default one generated by OpenNAS
			--U_BPF_0
			config_mem(0)  <= x"0002";
			config_mem(1)  <= x"700A";
			config_mem(2)  <= x"700A";
			config_mem(3)  <= x"2025";
			--U_BPF_1
			config_mem(4)  <= x"0003";
			config_mem(5)  <= x"6DDD";
			config_mem(6)  <= x"6DDD";
			config_mem(7)  <= x"2025";
			--U_BPF_2
			config_mem(8)  <= x"0002";
			config_mem(9)  <= x"7932";
			config_mem(10) <= x"7932";
			config_mem(11) <= x"2025";
			--U_BPF_3
			config_mem(12) <= x"0003";
			config_mem(13) <= x"76D8";
			config_mem(14) <= x"76D8";
			config_mem(15) <= x"2025";
			--U_BPF_4
			config_mem(16) <= x"0004";
			config_mem(17) <= x"6D40";
			config_mem(18) <= x"6D40";
			config_mem(19) <= x"2025";
			--U_BPF_5
			config_mem(20) <= x"0002";
			config_mem(21) <= x"606A";
			config_mem(22) <= x"606A";
			config_mem(23) <= x"2025";
			--U_BPF_6
			config_mem(24) <= x"0004";
			config_mem(25) <= x"762E";
			config_mem(26) <= x"762E";
			config_mem(27) <= x"2025";
			--U_BPF_7
			config_mem(28) <= x"0002";
			config_mem(29) <= x"684C";
			config_mem(30) <= x"684C";
			config_mem(31) <= x"2025";
			--U_BPF_8
			config_mem(32) <= x"0004";
			config_mem(33) <= x"7FD7";
			config_mem(34) <= x"7FD7";
			config_mem(35) <= x"2025";

		elsif rising_edge(clock) then
			if config_wren = '1' then
				for c_idx in 0 to CONFIG_OFFSET loop
					if to_integer(unsigned(config_addr)) = CONFIG_ADDRESS + c_idx then
						config_mem(c_idx) <= config_data;
					end if;
				end loop;
			end if;
		end if;
	end process;

	--Ideal cutoff: 36279,8110Hz - Real cutoff: 36278,4233Hz - Error: 0,0038%
	U_BPF_0 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 7,
			SAT => 63
		)
		Port Map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(0)(7 downto 0),
			spikes_div_fb   => config_mem(1),
			spikes_div_out  => config_mem(2),
			spikes_div_bpf  => config_mem(3),
			spike_in_slpf_p => spikes_in(1),
			spike_in_slpf_n => spikes_in(0),
			spike_in_shf_p  => '0',
			spike_in_shf_n  => '0',
			spike_out_p     => open,
			spike_out_n     => open,
			spike_out_lpf_p => lpf_spikes_0(1),
			spike_out_lpf_n => lpf_spikes_0(0)
		);

	--Ideal cutoff: 13340,7531Hz - Real cutoff: 13340,2132Hz - Error: 0,0040%
	U_BPF_1 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 8,
			SAT => 127
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(4)(7 downto 0),
			spikes_div_fb   => config_mem(5),
			spikes_div_out  => config_mem(6),
			spikes_div_bpf  => config_mem(7),
			spike_in_slpf_p => lpf_spikes_0(1),
			spike_in_slpf_n => lpf_spikes_0(0),
			spike_in_shf_p  => lpf_spikes_0(1),
			spike_in_shf_n  => lpf_spikes_0(0),
			spike_out_p     => spikes_out(1),
			spike_out_n     => spikes_out(0),
			spike_out_lpf_p => lpf_spikes_1(1),
			spike_out_lpf_n => lpf_spikes_1(0)
		);

	--Ideal cutoff: 4905,6400Hz - Real cutoff: 4905,4039Hz - Error: 0,0048%
	U_BPF_2 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 10,
			SAT => 511
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(8)(7 downto 0),
			spikes_div_fb   => config_mem(9),
			spikes_div_out  => config_mem(10),
			spikes_div_bpf  => config_mem(11),
			spike_in_slpf_p => lpf_spikes_1(1),
			spike_in_slpf_n => lpf_spikes_1(0),
			spike_in_shf_p  => lpf_spikes_1(1),
			spike_in_shf_n  => lpf_spikes_1(0),
			spike_out_p     => spikes_out(3),
			spike_out_n     => spikes_out(2),
			spike_out_lpf_p => lpf_spikes_2(1),
			spike_out_lpf_n => lpf_spikes_2(0)
		);

	--Ideal cutoff: 1803,8940Hz - Real cutoff: 1803,8340Hz - Error: 0,0033%
	U_BPF_3 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 11,
			SAT => 1023
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(12)(7 downto 0),
			spikes_div_fb   => config_mem(13),
			spikes_div_out  => config_mem(14),
			spikes_div_bpf  => config_mem(15),
			spike_in_slpf_p => lpf_spikes_2(1),
			spike_in_slpf_n => lpf_spikes_2(0),
			spike_in_shf_p  => lpf_spikes_2(1),
			spike_in_shf_n  => lpf_spikes_2(0),
			spike_out_p     => spikes_out(5),
			spike_out_n     => spikes_out(4),
			spike_out_lpf_p => lpf_spikes_3(1),
			spike_out_lpf_n => lpf_spikes_3(0)
		);

	--Ideal cutoff: 663,3250Hz - Real cutoff: 663,2873Hz - Error: 0,0057%
	U_BPF_4 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 12,
			SAT => 2047
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(16)(7 downto 0),
			spikes_div_fb   => config_mem(17),
			spikes_div_out  => config_mem(18),
			spikes_div_bpf  => config_mem(19),
			spike_in_slpf_p => lpf_spikes_3(1),
			spike_in_slpf_n => lpf_spikes_3(0),
			spike_in_shf_p  => lpf_spikes_3(1),
			spike_in_shf_n  => lpf_spikes_3(0),
			spike_out_p     => spikes_out(7),
			spike_out_n     => spikes_out(6),
			spike_out_lpf_p => lpf_spikes_4(1),
			spike_out_lpf_n => lpf_spikes_4(0)
		);

	--Ideal cutoff: 243,9168Hz - Real cutoff: 243,8986Hz - Error: 0,0074%
	U_BPF_5 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 14,
			SAT => 8191
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(20)(7 downto 0),
			spikes_div_fb   => config_mem(21),
			spikes_div_out  => config_mem(22),
			spikes_div_bpf  => config_mem(23),
			spike_in_slpf_p => lpf_spikes_4(1),
			spike_in_slpf_n => lpf_spikes_4(0),
			spike_in_shf_p  => lpf_spikes_4(1),
			spike_in_shf_n  => lpf_spikes_4(0),
			spike_out_p     => spikes_out(9),
			spike_out_n     => spikes_out(8),
			spike_out_lpf_p => lpf_spikes_5(1),
			spike_out_lpf_n => lpf_spikes_5(0)
		);

	--Ideal cutoff: 89,6927Hz - Real cutoff: 89,6877Hz - Error: 0,0055%
	U_BPF_6 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 15,
			SAT => 16383
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(24)(7 downto 0),
			spikes_div_fb   => config_mem(25),
			spikes_div_out  => config_mem(26),
			spikes_div_bpf  => config_mem(27),
			spike_in_slpf_p => lpf_spikes_5(1),
			spike_in_slpf_n => lpf_spikes_5(0),
			spike_in_shf_p  => lpf_spikes_5(1),
			spike_in_shf_n  => lpf_spikes_5(0),
			spike_out_p     => spikes_out(11),
			spike_out_n     => spikes_out(10),
			spike_out_lpf_p => lpf_spikes_6(1),
			spike_out_lpf_n => lpf_spikes_6(0)
		);

	--Ideal cutoff: 32,9816Hz - Real cutoff: 32,9800Hz - Error: 0,0051%
	U_BPF_7 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 17,
			SAT => 65535
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(28)(7 downto 0),
			spikes_div_fb   => config_mem(29),
			spikes_div_out  => config_mem(30),
			spikes_div_bpf  => config_mem(31),
			spike_in_slpf_p => lpf_spikes_6(1),
			spike_in_slpf_n => lpf_spikes_6(0),
			spike_in_shf_p  => lpf_spikes_6(1),
			spike_in_shf_n  => lpf_spikes_6(0),
			spike_out_p     => spikes_out(13),
			spike_out_n     => spikes_out(12),
			spike_out_lpf_p => lpf_spikes_7(1),
			spike_out_lpf_n => lpf_spikes_7(0)
		);

	--Ideal cutoff: 12,1280Hz - Real cutoff: 12,1274Hz - Error: 0,0049%
	U_BPF_8 : entity work.spikes_2BPF_fullGain
		Generic Map(
			GL  => 18,
			SAT => 131071
		)
		Port map(
			clk             => clock,
			rst             => not_rst,
			freq_div        => config_mem(32)(7 downto 0),
			spikes_div_fb   => config_mem(33),
			spikes_div_out  => config_mem(34),
			spikes_div_bpf  => config_mem(35),
			spike_in_slpf_p => lpf_spikes_7(1),
			spike_in_slpf_n => lpf_spikes_7(0),
			spike_in_shf_p  => lpf_spikes_7(1),
			spike_in_shf_n  => lpf_spikes_7(0),
			spike_out_p     => spikes_out(15),
			spike_out_n     => spikes_out(14),
			spike_out_lpf_p => lpf_spikes_8(1),
			spike_out_lpf_n => lpf_spikes_8(0)
		);

end CFBank_arq;
