
package OpenNas_top_pkg is
	constant CONFIG_BUS_BIT_WIDTH : integer := 16;
	constant AER_DATA_BUS_BIT_WIDTH : integer := 16;
	constant SPIKE_BUS_BIT_WIDTH : integer := 2;
end package OpenNas_top_pkg;

package body OpenNas_top_pkg is
	
end package body OpenNas_top_pkg;
