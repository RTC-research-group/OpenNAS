--/////////////////////////////////////////////////////////////////////////////////
--//                                                                             //
--//    Copyright � 2016  �ngel Francisco Jim�nez-Fern�ndez                      //
--//                                                                             //
--//    This file is part of OpenNAS.                                            //
--//                                                                             //
--//    OpenNAS is free software: you can redistribute it and/or modify          //
--//    it under the terms of the GNU General Public License as published by     //
--//    the Free Software Foundation, either version 3 of the License, or        //
--//    (at your option) any later version.                                      //
--//                                                                             //
--//    OpenNAS is distributed in the hope that it will be useful,               //
--//    but WITHOUT ANY WARRANTY; without even the implied warranty of           //
--//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.See the              //
--//    GNU General Public License for more details.                             //
--//                                                                             //
--//    You should have received a copy of the GNU General Public License        //
--//    along with OpenNAS. If not, see <http://www.gnu.org/licenses/>.          //
--//                                                                             //
--/////////////////////////////////////////////////////////////////////////////////

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity spikes_LPF_fullGain is
	Generic (
		GL             : INTEGER := 16; 
		SAT            : INTEGER := 32536
	);
    Port ( 
		clk            : in  STD_LOGIC;
		rst_n            : in  STD_LOGIC;
		freq_div       : in  STD_LOGIC_VECTOR(7 downto 0);
		spikes_div_fb  : in  STD_LOGIC_VECTOR(15 downto 0);
		spikes_div_out : in  STD_LOGIC_VECTOR(15 downto 0);
		spike_in_p     : in  STD_LOGIC;
		spike_in_n     : in  STD_LOGIC;
		spike_out_p    : out STD_LOGIC;
		spike_out_n    : out STD_LOGIC
	);
end spikes_LPF_fullGain;

architecture Behavioral of spikes_LPF_fullGain is
	
	signal int_spikes_p     : STD_LOGIC;
	signal int_spikes_n     : STD_LOGIC;
	signal spikes_out_tmp_p : STD_LOGIC;
	signal spikes_out_tmp_n : STD_LOGIC;
	signal spikes_fb_div_p  : STD_LOGIC;
	signal spikes_fb_div_n  : STD_LOGIC;

	begin

		U_OUT_DIV_out: entity work.spikes_div_BW
		Port Map (
			clk         => clk,
			rst_n         => rst_n,
			spikes_div  => spikes_div_out,
			spike_in_p  => spikes_out_tmp_p,
			spike_in_n  => spikes_out_tmp_n,
			spike_out_p => spike_out_p,
			spike_out_n => spike_out_n
		);

		U_FB_DIV: entity work.spikes_div_BW
		Port Map (
			clk         => clk,
			rst_n         => rst_n,
			spikes_div  => spikes_div_fb,
			spike_in_p  => spikes_out_tmp_p,
			spike_in_n  => spikes_out_tmp_n,
			spike_out_p => spikes_fb_div_p,
			spike_out_n => spikes_fb_div_n
		);

		U_DIF: entity work.AER_DIF
		Port Map (
			clk          =>clk,
			rst_n          =>rst_n,
			spkies_in_up =>spike_in_p,
			spikes_in_un =>spike_in_n,
			spikes_in_yp =>spikes_fb_div_p, 
			spikes_in_yn =>spikes_fb_div_n, 
			spikes_out_p =>int_spikes_p,
			spikes_out_n =>int_spikes_n
		);			  

		U_INT: entity work.Spike_Int_n_Gen_BW 
		Generic Map(
			GL          => GL, 
			SAT         => SAT
		)
		Port Map ( 
			clk         => clk,
			rst_n         => rst_n,
			freq_div    => freq_div,
			spike_in_p  => int_spikes_p,
			spike_in_n  => int_spikes_n,
			spike_out_p => spikes_out_tmp_p,
			spike_out_n => spikes_out_tmp_n
		);

end Behavioral;

