--/////////////////////////////////////////////////////////////////////////////////
--//                                                                             //
--//    Copyright � 2016  �ngel Francisco Jim�nez-Fern�ndez                      //
--//                                                                             //
--//    This file is part of OpenNAS.                                            //
--//                                                                             //
--//    OpenNAS is free software: you can redistribute it and/or modify          //
--//    it under the terms of the GNU General Public License as published by     //
--//    the Free Software Foundation, either version 3 of the License, or        //
--//    (at your option) any later version.                                      //
--//                                                                             //
--//    OpenNAS is distributed in the hope that it will be useful,               //
--//    but WITHOUT ANY WARRANTY; without even the implied warranty of           //
--//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.See the              //
--//    GNU General Public License for more details.                             //
--//                                                                             //
--//    You should have received a copy of the GNU General Public License        //
--//    along with OpenNAS. If not, see <http://www.gnu.org/licenses/>.          //
--//                                                                             //
--/////////////////////////////////////////////////////////////////////////////////

----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:34:54 02/24/2016 
-- Design Name: 
-- Module Name:    PDM2Spikes - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use work.OpenNas_top_pkg.all;
USE ieee.numeric_std.all;

entity PDM2Spikes is
	Generic (
		CONFIG_ADDRESS : integer := 16#0000#;
		CONFIG_OFFSET  : integer := 3;  -- Don't change this value
		SLPF_GL        : integer := 11;
		SLPF_SAT       : integer := 1023;
		SHPF_GL        : integer := 17;
		SHPF_SAT       : integer := 65535
	);
	Port (
		clk         : in  std_logic;
		rst_n         : in  std_logic;
		--PDM interface
		clock_div   : in  std_logic_vector(7 downto 0);
		pdm_clk     : out std_logic;
		pdm_dat     : in  std_logic;
		--Config Bus
		config_data : in  std_logic_vector(CONFIG_BUS_BIT_WIDTH - 1 downto 0);
		config_addr : in  std_logic_vector(CONFIG_BUS_BIT_WIDTH - 1 downto 0);
		config_wren : in  std_logic;
		--Output
		spikes_out  : out std_logic_vector(1 downto 0)
	);
end PDM2Spikes;

architecture Behavioral of PDM2Spikes is

	signal spikes_pdm      : std_logic_vector(1 downto 0);
	signal spikes_hpf_int  : std_logic_vector(1 downto 0);
	signal spikes_hpf_int2 : std_logic_vector(1 downto 0);
	signal spikes_int      : std_logic_vector(1 downto 0);
	--signal n_rst           : STD_LOGIC;

	-- Configurable signals
	type register_bank is array (0 to CONFIG_OFFSET) of std_logic_vector(CONFIG_BUS_BIT_WIDTH - 1 downto 0);
	signal config_mem : register_bank;
	
	begin

	--	n_rst <= not rst_n;
		
		U_Config_registers : process(clk, rst_n)
		begin
			if (rst_n = '0') then           -- In reset mode the parameter are the default one generated by OpenNAS
				for c_idx in 0 to (CONFIG_OFFSET) loop
					config_mem(c_idx) <= std_logic_vector(to_unsigned(PDM2Spikes_DEFAULT_parameter(c_idx), CONFIG_BUS_BIT_WIDTH));
				end loop;
	
			elsif rising_edge(clk) then
				if config_wren = '1' then
					for c_idx in 0 to CONFIG_OFFSET loop
						if to_integer(unsigned(config_addr)) = CONFIG_ADDRESS + c_idx then
							config_mem(c_idx) <= config_data;
						end if;
					end loop;
				end if;
			end if;
		end process;

		U_PDM_Interface: entity work.PDM_Interface
		Port Map (
			clk        => clk,
			rst_n        => rst_n,
			clock_div  => clock_div,
			pdm_clk    => pdm_clk,	
			pdm_dat    => pdm_dat,	
			spikes_out => spikes_pdm
		);

		U_SHPF1: entity work.Spikes_HPF
		Generic Map (
			GL          => SHPF_GL, 
			SAT         => SHPF_SAT
		)
		Port Map ( 
			clk         => clk,
			rst_n         => rst_n,
			freq_div    => config_mem(0)(7 downto 0),
			spike_in_p  => spikes_pdm(1),
			spike_in_n  => spikes_pdm(0),
			spike_out_p => spikes_hpf_int(1),
			spike_out_n => spikes_hpf_int(0)
		);

		U_SHPF2: entity work.Spikes_HPF
		Generic Map (
			GL          => SHPF_GL, 
			SAT         => SHPF_SAT
		)
		Port Map ( 
			clk         => clk,
			rst_n         => rst_n,
			freq_div    => config_mem(0)(7 downto 0),
			spike_in_p  => spikes_hpf_int(1),
			spike_in_n  => spikes_hpf_int(0),
			spike_out_p => spikes_hpf_int2(1),
			spike_out_n => spikes_hpf_int2(0)
		);
			
		U_LPF1: entity work.Spikes_2LPF_FullGain
		generic Map (
			GL             => SLPF_GL, 
			SAT            => SLPF_SAT
		)
		Port Map ( 
			clk            => clk,
			rst_n            => rst_n,
			freq_div       => config_mem(1)(7 downto 0),
			spikes_div_fb  => config_mem(2),
			spikes_div_out => config_mem(3),
			spike_in_p     => spikes_hpf_int2(1),
			spike_in_n     => spikes_hpf_int2(0),
			spike_out_p    => spikes_int(1),
			spike_out_n    => spikes_int(0)
		);

		spikes_out <= spikes_int;

end Behavioral;